// Placeholder for user_project_wrapper - no cambios aquí si estás usando TinyTapeout
module user_project_wrapper ();
endmodule
